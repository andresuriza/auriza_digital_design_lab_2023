module contador_manual_tb;
	reg dec;
	reg inc;
	reg reset;
	reg clk;
	wire [5:0] out;
	
	contador_regresivo modulo (.clk(clk),
					           .reset(reset),
								  .dec(dec),
								  .inc(inc),
					           .out(out));
								  
  initial begin
  dec = 0;
  dec = 1;
  #40
  dec = 0;
  dec = 1;
  #40
  dec = 0;
  dec = 1;
  #40
  dec = 0;
  dec = 1;
  #40
  inc = 0;
  inc = 1;
  #40
  inc = 0;
  inc = 1;
  
  end
 
 endmodule