module PosicionarBarcos #(parameter WIDTH = 4)(

input logic [WIDTH - 1:0] BarcosPersonasCoords,
input logic [WIDTH - 1:0] BarcosPCCoords,
input logic [2:0] DisparoCoords,

);





