module SeleccionarBarcos #(parameter WIDTH = 4)(

input logic [WIDTH - 1:0] NumBarcos
output logic [WIDTH - 1:0] NumBarcosTotal

);

4'b0000: NumBarcos = NumBarcosTotal

