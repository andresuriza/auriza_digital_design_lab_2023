module Jugando(input logic x,
					output logic jgdr, pc)
					
